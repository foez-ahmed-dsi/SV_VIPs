module test;
    initial begin
        $display("Testing");
    end
endmodule

